module rightAr_A_B(rightAr_R,A,B);

output [31:0] rightAr_R;
input [31:0] A,B;

wire Bfiveto31;

wire [31:0] conMux0,conMux1,conMux2,conMux3,conMux4;


two_to_one_mux mux0_1(conMux0[0],A[0],A[1],B[0]);
two_to_one_mux mux0_2(conMux0[1],A[1],A[2],B[0]);
two_to_one_mux mux0_3(conMux0[2],A[2],A[3],B[0]);
two_to_one_mux mux0_4(conMux0[3],A[3],A[4],B[0]);
two_to_one_mux mux0_5(conMux0[4],A[4],A[5],B[0]);
two_to_one_mux mux0_6(conMux0[5],A[5],A[6],B[0]);
two_to_one_mux mux0_7(conMux0[6],A[6],A[7],B[0]);
two_to_one_mux mux0_8(conMux0[7],A[7],A[8],B[0]);
two_to_one_mux mux0_9(conMux0[8],A[8],A[9],B[0]);
two_to_one_mux mux0_10(conMux0[9],A[9],A[10],B[0]);
two_to_one_mux mux0_11(conMux0[10],A[10],A[11],B[0]);
two_to_one_mux mux0_12(conMux0[11],A[11],A[12],B[0]);
two_to_one_mux mux0_13(conMux0[12],A[12],A[13],B[0]);
two_to_one_mux mux0_14(conMux0[13],A[13],A[14],B[0]);
two_to_one_mux mux0_15(conMux0[14],A[14],A[15],B[0]);
two_to_one_mux mux0_16(conMux0[15],A[15],A[16],B[0]);
two_to_one_mux mux0_17(conMux0[16],A[16],A[17],B[0]);
two_to_one_mux mux0_18(conMux0[17],A[17],A[18],B[0]);
two_to_one_mux mux0_19(conMux0[18],A[18],A[19],B[0]);
two_to_one_mux mux0_20(conMux0[19],A[19],A[20],B[0]);
two_to_one_mux mux0_21(conMux0[20],A[20],A[21],B[0]);
two_to_one_mux mux0_22(conMux0[21],A[21],A[22],B[0]);
two_to_one_mux mux0_23(conMux0[22],A[22],A[23],B[0]);
two_to_one_mux mux0_24(conMux0[23],A[23],A[24],B[0]);
two_to_one_mux mux0_25(conMux0[24],A[24],A[25],B[0]);
two_to_one_mux mux0_26(conMux0[25],A[25],A[26],B[0]);
two_to_one_mux mux0_27(conMux0[26],A[26],A[27],B[0]);
two_to_one_mux mux0_28(conMux0[27],A[27],A[28],B[0]);
two_to_one_mux mux0_29(conMux0[28],A[28],A[29],B[0]);
two_to_one_mux mux0_30(conMux0[29],A[29],A[30],B[0]);
two_to_one_mux mux0_31(conMux0[30],A[30],A[31],B[0]);
two_to_one_mux mux0_32(conMux0[31],A[31],A[31],B[0]);
					
two_to_one_mux mux1_1(conMux1[0],conMux0[0],conMux0[2],B[1]);
two_to_one_mux mux1_2(conMux1[1],conMux0[1],conMux0[3],B[1]);
two_to_one_mux mux1_3(conMux1[2],conMux0[2],conMux0[4],B[1]);
two_to_one_mux mux1_4(conMux1[3],conMux0[3],conMux0[5],B[1]);
two_to_one_mux mux1_5(conMux1[4],conMux0[4],conMux0[6],B[1]);
two_to_one_mux mux1_6(conMux1[5],conMux0[5],conMux0[7],B[1]);
two_to_one_mux mux1_7(conMux1[6],conMux0[6],conMux0[8],B[1]);
two_to_one_mux mux1_8(conMux1[7],conMux0[7],conMux0[9],B[1]);
two_to_one_mux mux1_9(conMux1[8],conMux0[8],conMux0[10],B[1]);
two_to_one_mux mux1_10(conMux1[9],conMux0[9],conMux0[11],B[1]);
two_to_one_mux mux1_11(conMux1[10],conMux0[10],conMux0[12],B[1]);
two_to_one_mux mux1_12(conMux1[11],conMux0[11],conMux0[13],B[1]);
two_to_one_mux mux1_13(conMux1[12],conMux0[12],conMux0[14],B[1]);
two_to_one_mux mux1_14(conMux1[13],conMux0[13],conMux0[15],B[1]);
two_to_one_mux mux1_15(conMux1[14],conMux0[14],conMux0[16],B[1]);
two_to_one_mux mux1_16(conMux1[15],conMux0[15],conMux0[17],B[1]);
two_to_one_mux mux1_17(conMux1[16],conMux0[16],conMux0[18],B[1]);
two_to_one_mux mux1_18(conMux1[17],conMux0[17],conMux0[19],B[1]);
two_to_one_mux mux1_19(conMux1[18],conMux0[18],conMux0[20],B[1]);
two_to_one_mux mux1_20(conMux1[19],conMux0[19],conMux0[21],B[1]);
two_to_one_mux mux1_21(conMux1[20],conMux0[20],conMux0[22],B[1]);
two_to_one_mux mux1_22(conMux1[21],conMux0[21],conMux0[23],B[1]);
two_to_one_mux mux1_23(conMux1[22],conMux0[22],conMux0[24],B[1]);
two_to_one_mux mux1_24(conMux1[23],conMux0[23],conMux0[25],B[1]);
two_to_one_mux mux1_25(conMux1[24],conMux0[24],conMux0[26],B[1]);
two_to_one_mux mux1_26(conMux1[25],conMux0[25],conMux0[27],B[1]);
two_to_one_mux mux1_27(conMux1[26],conMux0[26],conMux0[28],B[1]);
two_to_one_mux mux1_28(conMux1[27],conMux0[27],conMux0[29],B[1]);
two_to_one_mux mux1_29(conMux1[28],conMux0[28],conMux0[30],B[1]);
two_to_one_mux mux1_30(conMux1[29],conMux0[29],conMux0[31],B[1]);
two_to_one_mux mux1_31(conMux1[30],conMux0[30],conMux0[31],B[1]);
two_to_one_mux mux1_32(conMux1[31],conMux0[31],conMux0[31],B[1]);
					
two_to_one_mux mux2_1(conMux2[0],conMux1[0],conMux1[4],B[2]);
two_to_one_mux mux2_2(conMux2[1],conMux1[1],conMux1[5],B[2]);
two_to_one_mux mux2_3(conMux2[2],conMux1[2],conMux1[6],B[2]);
two_to_one_mux mux2_4(conMux2[3],conMux1[3],conMux1[7],B[2]);
two_to_one_mux mux2_5(conMux2[4],conMux1[4],conMux1[8],B[2]);
two_to_one_mux mux2_6(conMux2[5],conMux1[5],conMux1[9],B[2]);
two_to_one_mux mux2_7(conMux2[6],conMux1[6],conMux1[10],B[2]);
two_to_one_mux mux2_8(conMux2[7],conMux1[7],conMux1[11],B[2]);
two_to_one_mux mux2_9(conMux2[8],conMux1[8],conMux1[12],B[2]);
two_to_one_mux mux2_10(conMux2[9],conMux1[9],conMux1[13],B[2]);
two_to_one_mux mux2_11(conMux2[10],conMux1[10],conMux1[14],B[2]);
two_to_one_mux mux2_12(conMux2[11],conMux1[11],conMux1[15],B[2]);
two_to_one_mux mux2_13(conMux2[12],conMux1[12],conMux1[16],B[2]);
two_to_one_mux mux2_14(conMux2[13],conMux1[13],conMux1[17],B[2]);
two_to_one_mux mux2_15(conMux2[14],conMux1[14],conMux1[18],B[2]);
two_to_one_mux mux2_16(conMux2[15],conMux1[15],conMux1[19],B[2]);
two_to_one_mux mux2_17(conMux2[16],conMux1[16],conMux1[20],B[2]);
two_to_one_mux mux2_18(conMux2[17],conMux1[17],conMux1[21],B[2]);
two_to_one_mux mux2_19(conMux2[18],conMux1[18],conMux1[22],B[2]);
two_to_one_mux mux2_20(conMux2[19],conMux1[19],conMux1[23],B[2]);
two_to_one_mux mux2_21(conMux2[20],conMux1[20],conMux1[24],B[2]);
two_to_one_mux mux2_22(conMux2[21],conMux1[21],conMux1[25],B[2]);
two_to_one_mux mux2_23(conMux2[22],conMux1[22],conMux1[26],B[2]);
two_to_one_mux mux2_24(conMux2[23],conMux1[23],conMux1[27],B[2]);
two_to_one_mux mux2_25(conMux2[24],conMux1[24],conMux1[28],B[2]);
two_to_one_mux mux2_26(conMux2[25],conMux1[25],conMux1[29],B[2]);
two_to_one_mux mux2_27(conMux2[26],conMux1[26],conMux1[30],B[2]);
two_to_one_mux mux2_28(conMux2[27],conMux1[27],conMux1[31],B[2]);
two_to_one_mux mux2_29(conMux2[28],conMux1[28],conMux1[31],B[2]);
two_to_one_mux mux2_30(conMux2[29],conMux1[29],conMux1[31],B[2]);
two_to_one_mux mux2_31(conMux2[30],conMux1[30],conMux1[31],B[2]);
two_to_one_mux mux2_32(conMux2[31],conMux1[31],conMux1[31],B[2]);
				
two_to_one_mux mux3_1(conMux3[0],conMux2[0],conMux2[8],B[3]);
two_to_one_mux mux3_2(conMux3[1],conMux2[1],conMux2[9],B[3]);
two_to_one_mux mux3_3(conMux3[2],conMux2[2],conMux2[10],B[3]);
two_to_one_mux mux3_4(conMux3[3],conMux2[3],conMux2[11],B[3]);
two_to_one_mux mux3_5(conMux3[4],conMux2[4],conMux2[12],B[3]);
two_to_one_mux mux3_6(conMux3[5],conMux2[5],conMux2[13],B[3]);
two_to_one_mux mux3_7(conMux3[6],conMux2[6],conMux2[14],B[3]);
two_to_one_mux mux3_8(conMux3[7],conMux2[7],conMux2[15],B[3]);
two_to_one_mux mux3_9(conMux3[8],conMux2[8],conMux2[16],B[3]);
two_to_one_mux mux3_10(conMux3[9],conMux2[9],conMux2[17],B[3]);
two_to_one_mux mux3_11(conMux3[10],conMux2[10],conMux2[18],B[3]);
two_to_one_mux mux3_12(conMux3[11],conMux2[11],conMux2[19],B[3]);
two_to_one_mux mux3_13(conMux3[12],conMux2[12],conMux2[20],B[3]);
two_to_one_mux mux3_14(conMux3[13],conMux2[13],conMux2[21],B[3]);
two_to_one_mux mux3_15(conMux3[14],conMux2[14],conMux2[22],B[3]);
two_to_one_mux mux3_16(conMux3[15],conMux2[15],conMux2[23],B[3]);
two_to_one_mux mux3_17(conMux3[16],conMux2[16],conMux2[24],B[3]);
two_to_one_mux mux3_18(conMux3[17],conMux2[17],conMux2[25],B[3]);
two_to_one_mux mux3_19(conMux3[18],conMux2[18],conMux2[26],B[3]);
two_to_one_mux mux3_20(conMux3[19],conMux2[19],conMux2[27],B[3]);
two_to_one_mux mux3_21(conMux3[20],conMux2[20],conMux2[28],B[3]);
two_to_one_mux mux3_22(conMux3[21],conMux2[21],conMux2[29],B[3]);
two_to_one_mux mux3_23(conMux3[22],conMux2[22],conMux2[30],B[3]);
two_to_one_mux mux3_24(conMux3[23],conMux2[23],conMux2[31],B[3]);
two_to_one_mux mux3_25(conMux3[24],conMux2[24],conMux2[31],B[3]);
two_to_one_mux mux3_26(conMux3[25],conMux2[25],conMux2[31],B[3]);
two_to_one_mux mux3_27(conMux3[26],conMux2[26],conMux2[31],B[3]);
two_to_one_mux mux3_28(conMux3[27],conMux2[27],conMux2[31],B[3]);
two_to_one_mux mux3_29(conMux3[28],conMux2[28],conMux2[31],B[3]);
two_to_one_mux mux3_30(conMux3[29],conMux2[29],conMux2[31],B[3]);
two_to_one_mux mux3_31(conMux3[30],conMux2[30],conMux2[31],B[3]);
two_to_one_mux mux3_32(conMux3[31],conMux2[31],conMux2[31],B[3]);

two_to_one_mux mux4_1(conMux4[0],conMux3[0],conMux3[16],B[4]);
two_to_one_mux mux4_2(conMux4[1],conMux3[1],conMux3[17],B[4]);
two_to_one_mux mux4_3(conMux4[2],conMux3[2],conMux3[18],B[4]);
two_to_one_mux mux4_4(conMux4[3],conMux3[3],conMux3[19],B[4]);
two_to_one_mux mux4_5(conMux4[4],conMux3[4],conMux3[20],B[4]);
two_to_one_mux mux4_6(conMux4[5],conMux3[5],conMux3[21],B[4]);
two_to_one_mux mux4_7(conMux4[6],conMux3[6],conMux3[22],B[4]);
two_to_one_mux mux4_8(conMux4[7],conMux3[7],conMux3[23],B[4]);
two_to_one_mux mux4_9(conMux4[8],conMux3[8],conMux3[24],B[4]);
two_to_one_mux mux4_10(conMux4[9],conMux3[9],conMux3[25],B[4]);
two_to_one_mux mux4_11(conMux4[10],conMux3[10],conMux3[26],B[4]);
two_to_one_mux mux4_12(conMux4[11],conMux3[11],conMux3[27],B[4]);
two_to_one_mux mux4_13(conMux4[12],conMux3[12],conMux3[28],B[4]);
two_to_one_mux mux4_14(conMux4[13],conMux3[13],conMux3[29],B[4]);
two_to_one_mux mux4_15(conMux4[14],conMux3[14],conMux3[30],B[4]);
two_to_one_mux mux4_16(conMux4[15],conMux3[15],conMux3[31],B[4]);
two_to_one_mux mux4_17(conMux4[16],conMux3[16],conMux3[31],B[4]);
two_to_one_mux mux4_18(conMux4[17],conMux3[17],conMux3[31],B[4]);
two_to_one_mux mux4_19(conMux4[18],conMux3[18],conMux3[31],B[4]);
two_to_one_mux mux4_20(conMux4[19],conMux3[19],conMux3[31],B[4]);
two_to_one_mux mux4_21(conMux4[20],conMux3[20],conMux3[31],B[4]);
two_to_one_mux mux4_22(conMux4[21],conMux3[21],conMux3[31],B[4]);
two_to_one_mux mux4_23(conMux4[22],conMux3[22],conMux3[31],B[4]);
two_to_one_mux mux4_24(conMux4[23],conMux3[23],conMux3[31],B[4]);
two_to_one_mux mux4_25(conMux4[24],conMux3[24],conMux3[31],B[4]);
two_to_one_mux mux4_26(conMux4[25],conMux3[25],conMux3[31],B[4]);
two_to_one_mux mux4_27(conMux4[26],conMux3[26],conMux3[31],B[4]);
two_to_one_mux mux4_28(conMux4[27],conMux3[27],conMux3[31],B[4]);
two_to_one_mux mux4_29(conMux4[28],conMux3[28],conMux3[31],B[4]);
two_to_one_mux mux4_30(conMux4[29],conMux3[29],conMux3[31],B[4]);
two_to_one_mux mux4_31(conMux4[30],conMux3[30],conMux3[31],B[4]);
two_to_one_mux mux4_32(conMux4[31],conMux3[31],conMux3[31],B[4]);

or zeroALL(Bfiveto31,B[5],B[6],B[7],B[8],B[9],B[10],B[11],B[12],B[13],
			  B[14],B[15],B[16],B[17],B[18],B[19],B[20],B[21],B[22],B[23],B[24],
			  B[25],B[26],B[27],B[28],B[29],B[30],B[31]);

two_to_one_mux result1(rightAr_R[0],conMux4[0],0,Bfiveto31);
two_to_one_mux result2(rightAr_R[1],conMux4[1],0,Bfiveto31);
two_to_one_mux result3(rightAr_R[2],conMux4[2],0,Bfiveto31);
two_to_one_mux result4(rightAr_R[3],conMux4[3],0,Bfiveto31);
two_to_one_mux result5(rightAr_R[4],conMux4[4],0,Bfiveto31);
two_to_one_mux result6(rightAr_R[5],conMux4[5],0,Bfiveto31);
two_to_one_mux result7(rightAr_R[6],conMux4[6],0,Bfiveto31);
two_to_one_mux result8(rightAr_R[7],conMux4[7],0,Bfiveto31);
two_to_one_mux result9(rightAr_R[8],conMux4[8],0,Bfiveto31);
two_to_one_mux result10(rightAr_R[9],conMux4[9],0,Bfiveto31);
two_to_one_mux result11(rightAr_R[10],conMux4[10],0,Bfiveto31);
two_to_one_mux result12(rightAr_R[11],conMux4[11],0,Bfiveto31);
two_to_one_mux result13(rightAr_R[12],conMux4[12],0,Bfiveto31);
two_to_one_mux result14(rightAr_R[13],conMux4[13],0,Bfiveto31);
two_to_one_mux result15(rightAr_R[14],conMux4[14],0,Bfiveto31);
two_to_one_mux result16(rightAr_R[15],conMux4[15],0,Bfiveto31);
two_to_one_mux result17(rightAr_R[16],conMux4[16],0,Bfiveto31);
two_to_one_mux result18(rightAr_R[17],conMux4[17],0,Bfiveto31);
two_to_one_mux result19(rightAr_R[18],conMux4[18],0,Bfiveto31);
two_to_one_mux result20(rightAr_R[19],conMux4[19],0,Bfiveto31);
two_to_one_mux result21(rightAr_R[20],conMux4[20],0,Bfiveto31);
two_to_one_mux result22(rightAr_R[21],conMux4[21],0,Bfiveto31);
two_to_one_mux result23(rightAr_R[22],conMux4[22],0,Bfiveto31);
two_to_one_mux result24(rightAr_R[23],conMux4[23],0,Bfiveto31);
two_to_one_mux result25(rightAr_R[24],conMux4[24],0,Bfiveto31);
two_to_one_mux result26(rightAr_R[25],conMux4[25],0,Bfiveto31);
two_to_one_mux result27(rightAr_R[26],conMux4[26],0,Bfiveto31);
two_to_one_mux result28(rightAr_R[27],conMux4[27],0,Bfiveto31);
two_to_one_mux result29(rightAr_R[28],conMux4[28],0,Bfiveto31);
two_to_one_mux result30(rightAr_R[29],conMux4[29],0,Bfiveto31);
two_to_one_mux result31(rightAr_R[30],conMux4[30],0,Bfiveto31);
two_to_one_mux result32(rightAr_R[31],conMux4[31],0,Bfiveto31);


endmodule 