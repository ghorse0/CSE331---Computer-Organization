module or_A_B (or_A_B, A , B);

output [31:0] or_A_B ;
input [31:0] A,B ; 


or orOperation1(or_A_B[0],A[0],B[0]);
or orOperation2(or_A_B[1],A[1],B[1]);
or orOperation3(or_A_B[2],A[2],B[2]);
or orOperation4(or_A_B[3],A[3],B[3]);
or orOperation5(or_A_B[4],A[4],B[4]);
or orOperation6(or_A_B[5],A[5],B[5]);
or orOperation7(or_A_B[6],A[6],B[6]);
or orOperation8(or_A_B[7],A[7],B[7]);
or orOperation9(or_A_B[8],A[8],B[8]);
or orOperation10(or_A_B[9],A[9],B[9]);
or orOperation11(or_A_B[10],A[10],B[10]);
or orOperation12(or_A_B[11],A[11],B[11]);
or orOperation13(or_A_B[12],A[12],B[12]);
or orOperation14(or_A_B[13],A[13],B[13]);
or orOperation15(or_A_B[14],A[14],B[14]);
or orOperation16(or_A_B[15],A[15],B[15]);
or orOperation17(or_A_B[16],A[16],B[16]);
or orOperation18(or_A_B[17],A[17],B[17]);
or orOperation19(or_A_B[18],A[18],B[18]);
or orOperation20(or_A_B[19],A[19],B[19]);
or orOperation21(or_A_B[20],A[20],B[20]);
or orOperation22(or_A_B[21],A[21],B[21]);
or orOperation23(or_A_B[22],A[22],B[22]);
or orOperation24(or_A_B[23],A[23],B[23]);
or orOperation25(or_A_B[24],A[24],B[24]);
or orOperation26(or_A_B[25],A[25],B[25]);
or orOperation27(or_A_B[26],A[26],B[26]);
or orOperation28(or_A_B[27],A[27],B[27]);
or orOperation29(or_A_B[28],A[28],B[28]);
or orOperation30(or_A_B[29],A[29],B[29]);
or orOperation31(or_A_B[30],A[30],B[30]);
or orOperation32(or_A_B[31],A[31],B[31]);


endmodule 