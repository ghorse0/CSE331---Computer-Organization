module xor_A_B(xor_R , A , B);

output [31:0] xor_R;
input [31:0] A,B;


xor xorOperation1(xor_R[0],A[0],B[0]);
xor xorOperation2(xor_R[1],A[1],B[1]);
xor xorOperation3(xor_R[2],A[2],B[2]);
xor xorOperation4(xor_R[3],A[3],B[3]);
xor xorOperation5(xor_R[4],A[4],B[4]);
xor xorOperation6(xor_R[5],A[5],B[5]);
xor xorOperation7(xor_R[6],A[6],B[6]);
xor xorOperation8(xor_R[7],A[7],B[7]);
xor xorOperation9(xor_R[8],A[8],B[8]);
xor xorOperation10(xor_R[9],A[9],B[9]);
xor xorOperation11(xor_R[10],A[10],B[10]);
xor xorOperation12(xor_R[11],A[11],B[11]);
xor xorOperation13(xor_R[12],A[12],B[12]);
xor xorOperation14(xor_R[13],A[13],B[13]);
xor xorOperation15(xor_R[14],A[14],B[14]);
xor xorOperation16(xor_R[15],A[15],B[15]);
xor xorOperation17(xor_R[16],A[16],B[16]);
xor xorOperation18(xor_R[17],A[17],B[17]);
xor xorOperation19(xor_R[18],A[18],B[18]);
xor xorOperation20(xor_R[19],A[19],B[19]);
xor xorOperation21(xor_R[20],A[20],B[20]);
xor xorOperation22(xor_R[21],A[21],B[21]);
xor xorOperation23(xor_R[22],A[22],B[22]);
xor xorOperation24(xor_R[23],A[23],B[23]);
xor xorOperation25(xor_R[24],A[24],B[24]);
xor xorOperation26(xor_R[25],A[25],B[25]);
xor xorOperation27(xor_R[26],A[26],B[26]);
xor xorOperation28(xor_R[27],A[27],B[27]);
xor xorOperation29(xor_R[28],A[28],B[28]);
xor xorOperation30(xor_R[29],A[29],B[29]);
xor xorOperation31(xor_R[30],A[30],B[30]);
xor xorOperation32(xor_R[31],A[31],B[31]);



endmodule 