module nor_A_B(nor_R,A,B);

output [31:0] nor_R;
input [31:0] A,B;

nor norOperation1(nor_R[0],A[0],B[0]);
nor norOperation2(nor_R[1],A[1],B[1]);
nor norOperation3(nor_R[2],A[2],B[2]);
nor norOperation4(nor_R[3],A[3],B[3]);
nor norOperation5(nor_R[4],A[4],B[4]);
nor norOperation6(nor_R[5],A[5],B[5]);
nor norOperation7(nor_R[6],A[6],B[6]);
nor norOperation8(nor_R[7],A[7],B[7]);
nor norOperation9(nor_R[8],A[8],B[8]);
nor norOperation10(nor_R[9],A[9],B[9]);
nor norOperation11(nor_R[10],A[10],B[10]);
nor norOperation12(nor_R[11],A[11],B[11]);
nor norOperation13(nor_R[12],A[12],B[12]);
nor norOperation14(nor_R[13],A[13],B[13]);
nor norOperation15(nor_R[14],A[14],B[14]);
nor norOperation16(nor_R[15],A[15],B[15]);
nor norOperation17(nor_R[16],A[16],B[16]);
nor norOperation18(nor_R[17],A[17],B[17]);
nor norOperation19(nor_R[18],A[18],B[18]);
nor norOperation20(nor_R[19],A[19],B[19]);
nor norOperation21(nor_R[20],A[20],B[20]);
nor norOperation22(nor_R[21],A[21],B[21]);
nor norOperation23(nor_R[22],A[22],B[22]);
nor norOperation24(nor_R[23],A[23],B[23]);
nor norOperation25(nor_R[24],A[24],B[24]);
nor norOperation26(nor_R[25],A[25],B[25]);
nor norOperation27(nor_R[26],A[26],B[26]);
nor norOperation28(nor_R[27],A[27],B[27]);
nor norOperation29(nor_R[28],A[28],B[28]);
nor norOperation30(nor_R[29],A[29],B[29]);
nor norOperation31(nor_R[30],A[30],B[30]);
nor norOperation32(nor_R[31],A[31],B[31]);


endmodule 