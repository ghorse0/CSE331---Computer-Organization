module and_A_B (and_A_B, A , B);

output [31:0] and_A_B ;
input [31:0] A,B ; 


and andOperation1(and_A_B[0],A[0],B[0]);
and andOperation2(and_A_B[1],A[1],B[1]);
and andOperation3(and_A_B[2],A[2],B[2]);
and andOperation4(and_A_B[3],A[3],B[3]);
and andOperation5(and_A_B[4],A[4],B[4]);
and andOperation6(and_A_B[5],A[5],B[5]);
and andOperation7(and_A_B[6],A[6],B[6]);
and andOperation8(and_A_B[7],A[7],B[7]);
and andOperation9(and_A_B[8],A[8],B[8]);
and andOperation10(and_A_B[9],A[9],B[9]);
and andOperation11(and_A_B[10],A[10],B[10]);
and andOperation12(and_A_B[11],A[11],B[11]);
and andOperation13(and_A_B[12],A[12],B[12]);
and andOperation14(and_A_B[13],A[13],B[13]);
and andOperation15(and_A_B[14],A[14],B[14]);
and andOperation16(and_A_B[15],A[15],B[15]);
and andOperation17(and_A_B[16],A[16],B[16]);
and andOperation18(and_A_B[17],A[17],B[17]);
and andOperation19(and_A_B[18],A[18],B[18]);
and andOperation20(and_A_B[19],A[19],B[19]);
and andOperation21(and_A_B[20],A[20],B[20]);
and andOperation22(and_A_B[21],A[21],B[21]);
and andOperation23(and_A_B[22],A[22],B[22]);
and andOperation24(and_A_B[23],A[23],B[23]);
and andOperation25(and_A_B[24],A[24],B[24]);
and andOperation26(and_A_B[25],A[25],B[25]);
and andOperation27(and_A_B[26],A[26],B[26]);
and andOperation28(and_A_B[27],A[27],B[27]);
and andOperation29(and_A_B[28],A[28],B[28]);
and andOperation30(and_A_B[29],A[29],B[29]);
and andOperation31(and_A_B[30],A[30],B[30]);
and andOperation32(and_A_B[31],A[31],B[31]);


endmodule 